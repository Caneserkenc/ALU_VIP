package alu_pkg;

     import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "agent/alu_seq_item.svh"
    `include "sequence/alu_base_sequence.svh"

    `include "agent/alu_driver.svh"

    `include "agent/alu_monitor.svh"


    
    `include "agent/alu_agent.svh"
    `include "scoreboard/alu_scoreboard.svh"
    `include "env/alu_env.svh"

    `include "test/alu_test.svh"



endpackage